module idle_mem (
    input [3:0] step,
    input [7:0] ram_addr,
    output [0:15] ram_data [131:0]
);

    parameter [0:15] step0 [21384:0] = {
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00080, 16'd010C1, 16'd01102, 16'd01102, 16'd010C1, 16'd00080, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd01081, 16'd01081, 16'd01081, 16'd01041, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00080, 16'd010C1, 16'd01102, 16'd01102, 16'd010C1, 16'd00080, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd01081, 16'd01081, 16'd01081, 16'd01041, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00080, 16'd010C1, 16'd010C1, 16'd01101, 16'd010C1, 16'd00080, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd01081, 16'd01081, 16'd01081, 16'd01041, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00080, 16'd01081, 16'd010C1, 16'd010C1, 16'd010C1, 16'd00080, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd01081, 16'd01081, 16'd01081, 16'd01041, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00080, 16'd01081, 16'd01081, 16'd00081, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd01081, 16'd02081, 16'd02081, 16'd01041, 16'd01040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00080, 16'd00080, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd01040, 16'd01040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd01041, 16'd02081, 16'd02081, 16'd01041, 16'd01040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd01040, 16'd01080, 16'd01081, 16'd01080, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd01041, 16'd02081, 16'd02081, 16'd02041, 16'd01041, 16'd01040, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd01040, 16'd01081, 16'd02081, 16'd01081, 16'd01040, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd01041, 16'd02081, 16'd02081, 16'd02041, 16'd01041, 16'd01040, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd01041, 16'd02081, 16'd02081, 16'd02081, 16'd01041, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01040, 16'd01041, 16'd01041, 16'd01041, 16'd01041, 16'd01040, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01040, 16'd02081, 16'd02081, 16'd030C2, 16'd02081, 16'd01041, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01041, 16'd01041, 16'd01040, 16'd01040, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01040, 16'd02081, 16'd030C2, 16'd030C2, 16'd03082, 16'd02081, 16'd01040, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02040, 16'd02081, 16'd030C2, 16'd040C2, 16'd03082, 16'd02081, 16'd01040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02040, 16'd03081, 16'd040C2, 16'd040C2, 16'd03082, 16'd02081, 16'd01040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02040, 16'd03041, 16'd04082, 16'd040C2, 16'd03082, 16'd02081, 16'd01040, 16'd01000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02040, 16'd02041, 16'd03081, 16'd03081, 16'd03081, 16'd02041, 16'd02040, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02040, 16'd03041, 16'd03081, 16'd03041, 16'd02040, 16'd02040, 16'd01000, 16'd01000, 16'd02040, 16'd02041, 16'd02041, 16'd02041, 16'd02000, 16'd01000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02040, 16'd02040, 16'd02040, 16'd02040, 16'd02000, 16'd02000, 16'd02000, 16'd02040, 16'd03041, 16'd03041, 16'd03041, 16'd02041, 16'd01000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02040, 16'd02041, 16'd03041, 16'd03082, 16'd03042, 16'd02041, 16'd02000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02040, 16'd02041, 16'd03041, 16'd03082, 16'd03042, 16'd02041, 16'd02000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02040, 16'd02041, 16'd02041, 16'd02041, 16'd02041, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00080, 16'd00080, 16'd00080, 16'd00080,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00080, 16'd00080, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02041, 16'd02001, 16'd01000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00080, 16'd00080, 16'd00080, 16'd00080,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00081, 16'd00081, 16'd00080, 16'd00080, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00080, 16'd00080, 16'd00080, 16'd00080,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00081, 16'd000C1, 16'd000C1, 16'd000C1, 16'd00080, 16'd00080, 16'd00080, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00080, 16'd00080, 16'd00080, 16'd00080,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00081, 16'd000C1, 16'd000C1, 16'd000C1, 16'd00080, 16'd00080, 16'd00080, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00080, 16'd00080, 16'd00080, 16'd00080,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00080, 16'd00081, 16'd000C1, 16'd000C0, 16'd000C0, 16'd00080, 16'd00080, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00080, 16'd00080, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01040, 16'd01040, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00080, 16'd00080, 16'd00080, 16'd00080,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00080, 16'd00080, 16'd00080, 16'd000C0, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00080, 16'd00080, 16'd000C1, 16'd000C1, 16'd000C1, 16'd000C1, 16'd00081, 16'd01081, 16'd01081, 16'd01081, 16'd01081, 16'd01041, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01041, 16'd02041, 16'd02041, 16'd01041, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00040, 16'd00040, 16'd00040, 16'd00080, 16'd00080, 16'd000C1, 16'd00101, 16'd00102, 16'd00102, 16'd01102, 16'd01102, 16'd010C2, 16'd010C2, 16'd010C1, 16'd01081, 16'd01081, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd02041, 16'd02082, 16'd02082, 16'd02041, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd000C1, 16'd00101, 16'd00102, 16'd00142, 16'd00142, 16'd01142, 16'd01102, 16'd01102, 16'd01102, 16'd01102, 16'd010C1, 16'd01081, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd01040, 16'd02081, 16'd03082, 16'd03082, 16'd02081, 16'd01041, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd000C0, 16'd000C0, 16'd000C0, 16'd00101, 16'd00101, 16'd00102, 16'd00142, 16'd00142, 16'd01142, 16'd01102, 16'd01102, 16'd01102, 16'd01102, 16'd010C1, 16'd01081, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd01040, 16'd02081, 16'd02082, 16'd02082, 16'd02081, 16'd01041, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00080, 16'd00080, 16'd000C0, 16'd000C0, 16'd00100, 16'd00101, 16'd00101, 16'd00101, 16'd00101, 16'd00102, 16'd01102, 16'd01102, 16'd01102, 16'd01101, 16'd010C1, 16'd010C1, 16'd01081, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01041, 16'd02081, 16'd02081, 16'd02041, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd00000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00080, 16'd000C0, 16'd00100, 16'd00100, 16'd00101, 16'd00101, 16'd00101, 16'd00101, 16'd00101, 16'd00101, 16'd000C1, 16'd000C1, 16'd010C1, 16'd010C1, 16'd010C1, 16'd01081, 16'd00080, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01041, 16'd01041, 16'd01041, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00080, 16'd00100, 16'd00141, 16'd00181, 16'd00181, 16'd00141, 16'd00100, 16'd000C0, 16'd000C0, 16'd000C0, 16'd000C0, 16'd000C0, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd000C0, 16'd00140, 16'd001C2, 16'd00203, 16'd00244, 16'd00203, 16'd00182, 16'd00101, 16'd000C0, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00080, 16'd010C1, 16'd02142, 16'd021C3, 16'd03203, 16'd03203, 16'd03203, 16'd02203, 16'd02243, 16'd02285, 16'd02307, 16'd02388, 16'd02388, 16'd02307, 16'd01244, 16'd00141, 16'd000C0, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01081, 16'd031C4, 16'd062C8, 16'd093CB, 16'd0A48D, 16'd0A48D, 16'd0A48D, 16'd0948C, 16'd0948C, 16'd0950E, 16'd0A550, 16'd0A591, 16'd09590, 16'd0748C, 16'd04348, 16'd011C3, 16'd00100, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00040, 16'd00040, 16'd00040, 16'd00081, 16'd01081, 16'd010C2, 16'd01082, 16'd01041, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01102, 16'd062C8, 16'd0C4CF, 16'd11655, 16'd13758, 16'd14799, 16'd13798, 16'd12757, 16'd11757, 16'd127D8, 16'd1281A, 16'd1281A, 16'd11799, 16'd0D653, 16'd0844C, 16'd03285, 16'd00140, 16'd00080, 16'd00080, 16'd000C0, 16'd000C0, 16'd00080, 16'd00080, 16'd00040, 16'd00040, 16'd00080, 16'd010C1, 16'd02103, 16'd03144, 16'd03103, 16'd020C2, 16'd00041, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd02143, 16'd0A3CC, 16'd12696, 16'd1991F, 16'd1DA63, 16'd1DAA4, 16'd1CAA3, 16'd1AA62, 16'd1AA21, 16'd1AAA3, 16'd1BAA4, 16'd1BAA4, 16'd199E1, 16'd1381A, 16'd0B590, 16'd04307, 16'd00180, 16'd000C0, 16'd00080, 16'd000C0, 16'd000C0, 16'd000C0, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd02102, 16'd03144, 16'd04185, 16'd04185, 16'd03103, 16'd01081, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd03184, 16'd0C48F, 16'd1781C, 16'd20B27, 16'd25CED, 16'd25D2E, 16'd23CEC, 16'd21CAA, 16'd20C6A, 16'd21CAB, 16'd22CEC, 16'd22CAC, 16'd1FBA8, 16'd1895F, 16'd0F653, 16'd05388, 16'd00181, 16'd000C0, 16'd00080, 16'd000C0, 16'd00100, 16'd000C0, 16'd00080, 16'd00080, 16'd00080, 16'd010C1, 16'd02103, 16'd04185, 16'd05206, 16'd051C6, 16'd03144, 16'd01082, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd04184, 16'd0E511, 16'd1B920, 16'd25CAC, 16'd2AE73, 16'd2AEB4, 16'd28E72, 16'd25DEF, 16'd24DAE, 16'd25DF0, 16'd26E31, 16'd26DF0, 16'd23CED, 16'd1BA63, 16'd11716, 16'd063C9, 16'd00181, 16'd00080, 16'd00080, 16'd000C0, 16'd00100, 16'd000C0, 16'd000C0, 16'd00080, 16'd00080, 16'd010C1, 16'd02143, 16'd04185, 16'd05206, 16'd051C6, 16'd03144, 16'd020C2, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd041C5, 16'd10592, 16'd1D9E3, 16'd28DB0, 16'd2DF77, 16'd2DFB7, 16'd2AF34, 16'd26E71, 16'd25DF0, 16'd26E71, 16'd28EB3, 16'd29EB3, 16'd25D6F, 16'd1DAE4, 16'd12717, 16'd073C9, 16'd00180, 16'd00080, 16'd00080, 16'd000C0, 16'd00100, 16'd000C0, 16'd000C0, 16'd00080, 16'd00080, 16'd000C0, 16'd02102, 16'd03184, 16'd041C5, 16'd04185, 16'd03144, 16'd020C3, 16'd01081, 16'd01041, 16'd00041, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd01000, 16'd01000, 16'd01000, 16'd01000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd041C5, 16'd115D3, 16'd1FA64, 16'd2BE33, 16'd30FF9, 16'd2FFF9, 16'd2BF35, 16'd26E31, 16'd24DEF, 16'd26E71, 16'd28EB3, 16'd29EF4, 16'd27DB0, 16'd1EAE5, 16'd12757, 16'd07389, 16'd00140, 16'd00040, 16'd00040, 16'd000C0, 16'd00100, 16'd00100, 16'd000C0, 16'd000C0, 16'd00080, 16'd000C0, 16'd010C1, 16'd02102, 16'd03143, 16'd03143, 16'd03103, 16'd020C3, 16'd020C2, 16'd02082, 16'd01081, 16'd01040, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd01000, 16'd01000, 16'd01000, 16'd01000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd041C5, 16'd115D4, 16'd20AA6, 16'd2CE74, 16'd31FFA, 16'd30FF9, 16'd2BF35, 16'd25DF0, 16'd23DAE, 16'd25DF0, 16'd28EB3, 16'd2AEF4, 16'd27DB0, 16'd1EAE5, 16'd13717, 16'd07389, 16'd00100, 16'd00040, 16'd00040, 16'd000C0, 16'd00100, 16'd00100, 16'd00100, 16'd000C0, 16'd000C0, 16'd000C0, 16'd00080, 16'd01081, 16'd010C1, 16'd010C2, 16'd020C2, 16'd02103, 16'd03103, 16'd030C3, 16'd02082, 16'd01041, 16'd01000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd01000, 16'd01000, 16'd01000, 16'd01000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd041C5, 16'd12614, 16'd21AA6, 16'd2DEB5, 16'd32FFB, 16'd30FF9, 16'd2AEF4, 16'd25DAF, 16'd23D2D, 16'd24DAF, 16'd28E72, 16'd29EB4, 16'd27DB0, 16'd1EAE5, 16'd13717, 16'd07349, 16'd00100, 16'd00040, 16'd00040, 16'd000C0, 16'd00100, 16'd00100, 16'd00100, 16'd000C0, 16'd000C0, 16'd000C0, 16'd00080, 16'd00040, 16'd00040, 16'd00080, 16'd010C2, 16'd02103, 16'd03144, 16'd03103, 16'd030C3, 16'd02081, 16'd01000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd041C5, 16'd12614, 16'd21AA6, 16'd2DEB5, 16'd32FFB, 16'd30FF9, 16'd2BEF4, 16'd25DAF, 16'd23D2D, 16'd25DAF, 16'd28E72, 16'd29EB3, 16'd27DB0, 16'd1EAE5, 16'd13717, 16'd07389, 16'd00100, 16'd00040, 16'd00040, 16'd000C0, 16'd00100, 16'd00100, 16'd00100, 16'd00100, 16'd000C0, 16'd000C0, 16'd00080, 16'd00040, 16'd00040, 16'd00040, 16'd01081, 16'd02103, 16'd03144, 16'd03103, 16'd030C3, 16'd02081, 16'd01000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd041C5, 16'd125D4, 16'd21AA6, 16'd2DE74, 16'd32FFA, 16'd30FF9, 16'd2BEF4, 16'd26DAF, 16'd24D6D, 16'd25DAF, 16'd28E72, 16'd2AEB3, 16'd27DB0, 16'd1FAE6, 16'd13758, 16'd073CA, 16'd00141, 16'd00080, 16'd00080, 16'd000C0, 16'd00100, 16'd00100, 16'd00100, 16'd00100, 16'd00100, 16'd000C0, 16'd000C0, 16'd00080, 16'd00040, 16'd00080, 16'd01081, 16'd020C2, 16'd02103, 16'd03103, 16'd02082, 16'd01041, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd041C5, 16'd115D4, 16'd20A25, 16'd2CE33, 16'd31FB9, 16'd30FB8, 16'd2BEF4, 16'd27DF0, 16'd25D6E, 16'd26DF0, 16'd29E72, 16'd2AE73, 16'd27D6F, 16'd1EAE6, 16'd13758, 16'd0740B, 16'd001C2, 16'd000C1, 16'd00080, 16'd000C0, 16'd000C0, 16'd000C0, 16'd00100, 16'd00100, 16'd00101, 16'd00101, 16'd000C1, 16'd000C1, 16'd000C1, 16'd00081, 16'd01081, 16'd010C2, 16'd020C2, 16'd02082, 16'd01081, 16'd01040, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd041C5, 16'd10553, 16'd1E9E3, 16'd2AD70, 16'd2FF37, 16'd2FF77, 16'd2BEB3, 16'd27DB0, 16'd25D6E, 16'd27DB0, 16'd29E31, 16'd29E32, 16'd26D2E, 16'd1EAA5, 16'd12758, 16'd0744C, 16'd00204, 16'd00101, 16'd000C0, 16'd000C0, 16'd000C0, 16'd000C0, 16'd000C0, 16'd00101, 16'd00141, 16'd00141, 16'd00102, 16'd00102, 16'd01102, 16'd010C2, 16'd010C2, 16'd01081, 16'd01081, 16'd01041, 16'd01041, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd04184, 16'd0F511, 16'd1C920, 16'd27C6D, 16'd2CE33, 16'd2CE73, 16'd29DF1, 16'd26D2E, 16'd24CED, 16'd26D2E, 16'd27D6F, 16'd27D6F, 16'd24C6C, 16'd1CA23, 16'd11758, 16'd0644C, 16'd00245, 16'd00141, 16'd000C0, 16'd000C0, 16'd000C0, 16'd000C0, 16'd000C0, 16'd00101, 16'd00142, 16'd00142, 16'd00142, 16'd01142, 16'd01102, 16'd01102, 16'd010C2, 16'd00081, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd03144, 16'd0D48F, 16'd1981C, 16'd23B28, 16'd27CAD, 16'd27CEE, 16'd25C6C, 16'd22BE9, 16'd21BA8, 16'd22BE9, 16'd23C2A, 16'd23BEA, 16'd20B27, 16'd1991F, 16'd0F696, 16'd0640C, 16'd00245, 16'd00141, 16'd00100, 16'd000C0, 16'd00080, 16'd00080, 16'd000C0, 16'd00101, 16'd00102, 16'd00142, 16'd00142, 16'd01143, 16'd01143, 16'd01102, 16'd010C2, 16'd00041, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd02103, 16'd0A38C, 16'd14697, 16'd1B920, 16'd1FA64, 16'd1FAA5, 16'd1DA23, 16'd1B9E1, 16'd1B9A0, 16'd1B9A1, 16'd1C9E2, 16'd1C9A2, 16'd1A91F, 16'd14799, 16'd0C591, 16'd0438A, 16'd00204, 16'd00141, 16'd000C0, 16'd000C0, 16'd00080, 16'd00080, 16'd00080, 16'd000C1, 16'd00101, 16'd00101, 16'd00102, 16'd01102, 16'd01102, 16'd010C2, 16'd00081, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd020C2, 16'd072C9, 16'd0D4D0, 16'd13697, 16'd1579A, 16'd1579A, 16'd14759, 16'd13717, 16'd126D6, 16'd136D7, 16'd13717, 16'd13717, 16'd12696, 16'd0E591, 16'd0840C, 16'd032C7, 16'd001C3, 16'd00101, 16'd000C0, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd000C1, 16'd000C1, 16'd000C1, 16'd000C1, 16'd010C1, 16'd00081, 16'd00081, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01081, 16'd041C5, 16'd0730A, 16'd0A44D, 16'd0B4CF, 16'd0B4CF, 16'd0B44E, 16'd0A40C, 16'd0A40C, 16'd0A40C, 16'd0A44D, 16'd0A44D, 16'd0940C, 16'd0734A, 16'd04287, 16'd011C4, 16'd00141, 16'd000C0, 16'd00080, 16'd00080, 16'd00040, 16'd00040, 16'd00040, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00081, 16'd00081, 16'd00041, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd010C2, 16'd02184, 16'd03205, 16'd03246, 16'd03246, 16'd03205, 16'd031C4, 16'd031C3, 16'd031C3, 16'd031C4, 16'd031C4, 16'd031C4, 16'd02183, 16'd01142, 16'd00101, 16'd000C0, 16'd000C0, 16'd00080, 16'd00080, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00080, 16'd000C1, 16'd000C0, 16'd000C0, 16'd00080, 16'd00040, 16'd00040, 16'd00040, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00040, 16'd00040, 16'd01081, 16'd01081, 16'd01081, 16'd01040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd01081, 16'd010C1, 16'd020C2, 16'd020C2, 16'd01081, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00080, 16'd00080, 16'd00080, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd01081, 16'd020C2, 16'd02102, 16'd02102, 16'd020C1, 16'd01040, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd01081, 16'd02102, 16'd03103, 16'd02102, 16'd020C2, 16'd01041, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01040, 16'd01040, 16'd01040, 16'd01040, 16'd00040, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd01040, 16'd01081, 16'd010C1, 16'd020C2, 16'd02102, 16'd020C2, 16'd01081, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01040, 16'd02041, 16'd02081, 16'd03082, 16'd02081, 16'd01040, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd01040, 16'd01040, 16'd01081, 16'd02081, 16'd02081, 16'd020C1, 16'd020C2, 16'd020C1, 16'd01081, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01041, 16'd03082, 16'd040C3, 16'd040C3, 16'd030C2, 16'd02041, 16'd01040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01040, 16'd01040, 16'd02081, 16'd020C2, 16'd030C2, 16'd020C2, 16'd020C1, 16'd01081, 16'd01041, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd02081, 16'd040C2, 16'd05103, 16'd05104, 16'd040C3, 16'd03081, 16'd01040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01040, 16'd02080, 16'd020C1, 16'd030C2, 16'd03103, 16'd03102, 16'd020C1, 16'd01041, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd02081, 16'd040C3, 16'd05104, 16'd06144, 16'd04103, 16'd03081, 16'd01040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01040, 16'd02080, 16'd030C1, 16'd03102, 16'd04103, 16'd03102, 16'd02081, 16'd01040, 16'd00000, 16'd00040, 16'd00081, 16'd010C2, 16'd02103, 16'd02103, 16'd010C2, 16'd00081, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd02041, 16'd030C2, 16'd05103, 16'd05103, 16'd040C2, 16'd03081, 16'd02040, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01040, 16'd02081, 16'd030C2, 16'd03102, 16'd030C2, 16'd01081, 16'd00000, 16'd00000, 16'd01081, 16'd04144, 16'd07248, 16'd092CA, 16'd082C9, 16'd06207, 16'd03143, 16'd00080, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01041, 16'd03082, 16'd040C2, 16'd040C2, 16'd03082, 16'd03041, 16'd02040, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd01040, 16'd02041, 16'd02081, 16'd020C2, 16'd02081, 16'd01041, 16'd00000, 16'd00040, 16'd03103, 16'd08289, 16'd0E44F, 16'd12513, 16'd114D2, 16'd0C3CD, 16'd06206, 16'd010C1, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd02041, 16'd02041, 16'd03041, 16'd02041, 16'd02040, 16'd02040, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd01040, 16'd01041, 16'd01041, 16'd01041, 16'd00040, 16'd00000, 16'd00040, 16'd051C5, 16'd0D40E, 16'd16657, 16'd1C79D, 16'd1A75B, 16'd13554, 16'd0A2CA, 16'd020C2, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd02000, 16'd02040, 16'd02040, 16'd02040, 16'd02040, 16'd02040, 16'd02040, 16'd02040, 16'd02040, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00080, 16'd06247, 16'd12553, 16'd1D81E, 16'd249E5, 16'd22963, 16'd196DA, 16'd0D3CD, 16'd02102, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd02000, 16'd02040, 16'd02040, 16'd02040, 16'd02040, 16'd02040, 16'd02040, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00080, 16'd07288, 16'd15616, 16'd22963, 16'd2AB6B, 16'd28AE9, 16'd1D7DE, 16'd0F44F, 16'd03103, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd02040, 16'd02040, 16'd02040, 16'd02040, 16'd02000, 16'd02040, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00080, 16'd082C9, 16'd16657, 16'd25A26, 16'd2DC2F, 16'd2BBAC, 16'd1F8A0, 16'd10490, 16'd03143, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01040, 16'd01040, 16'd01040, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd082C9, 16'd17698, 16'd26A67, 16'd2ECB0, 16'd2CBEE, 16'd208E1, 16'd10491, 16'd03143, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01040, 16'd01040, 16'd01040, 16'd01040, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd01040, 16'd01040, 16'd01081, 16'd00080, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd08288, 16'd17698, 16'd26A67, 16'd2FCB0, 16'd2CC2E, 16'd208E2, 16'd104D1, 16'd03143, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01040, 16'd01040, 16'd01040, 16'd01040, 16'd01040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd01081, 16'd01081, 16'd01081, 16'd00080, 16'd00080, 16'd00080, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd08288, 16'd16657, 16'd25A67, 16'd2ECB0, 16'd2CC2E, 16'd208E1, 16'd104D1, 16'd03143, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01040, 16'd01040, 16'd01040, 16'd01040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd01081, 16'd010C1, 16'd010C1, 16'd000C1, 16'd00080, 16'd00080, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd07248, 16'd16657, 16'd25A67, 16'd2ECB0, 16'd2CC2E, 16'd208E1, 16'd104D1, 16'd03143, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd01040, 16'd01040, 16'd01040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00081, 16'd01081, 16'd010C1, 16'd000C1, 16'd000C1, 16'd000C0, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd07247, 16'd16657, 16'd24A26, 16'd2DCAF, 16'd2BBED, 16'd1F8E1, 16'd104D1, 16'd03143, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd01040, 16'd01040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00080, 16'd00080, 16'd00081, 16'd000C1, 16'd000C1, 16'd000C1, 16'd00080, 16'd00000, 16'd00000, 16'd00000, 16'd07247, 16'd15616, 16'd239E5, 16'd2CC2E, 16'd29BAC, 16'd1E8A0, 16'd0F490, 16'd03143, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00080, 16'd00081, 16'd000C1, 16'd000C1, 16'd00080, 16'd00000, 16'd00000, 16'd00040, 16'd07247, 16'd145D5, 16'd229A4, 16'd2ABED, 16'd28B2A, 16'd1D85F, 16'd0F490, 16'd03143, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00080, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00080, 16'd000C1, 16'd000C1, 16'd00080, 16'd00000, 16'd00000, 16'd00040, 16'd07247, 16'd135D5, 16'd20962, 16'd28B6B, 16'd26AE9, 16'd1C81E, 16'd0E44F, 16'd03143, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00080, 16'd00080, 16'd00080, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00080, 16'd000C1, 16'd00101, 16'd000C0, 16'd00000, 16'd00000, 16'd00040, 16'd06247, 16'd13594, 16'd20922, 16'd27B2A, 16'd25AA8, 16'd1B7DD, 16'd0E44F, 16'd03143, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00040, 16'd00040, 16'd00000, 16'd00040, 16'd00080, 16'd000C1, 16'd00101, 16'd000C0, 16'd00000, 16'd00000, 16'd00040, 16'd06247, 16'd13594, 16'd1F921, 16'd27B2A, 16'd25AA7, 16'd1B7DD, 16'd0E44F, 16'd03143, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd03000, 16'd03000, 16'd03000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00040, 16'd00000, 16'd00000, 16'd00040, 16'd00080, 16'd000C1, 16'd00101, 16'd000C0, 16'd00000, 16'd00000, 16'd00040, 16'd06247, 16'd12594, 16'd1F921, 16'd27B29, 16'd25A67, 16'd1B7DD, 16'd0E44F, 16'd03143, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd03000, 16'd03000, 16'd03000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00040, 16'd00000, 16'd00000, 16'd00040, 16'd00080, 16'd000C1, 16'd00101, 16'd000C0, 16'd00000, 16'd00000, 16'd00040, 16'd06247, 16'd12594, 16'd1F921, 16'd27B29, 16'd25A67, 16'd1B7DD, 16'd0E44F, 16'd03143, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd03000, 16'd03000, 16'd03000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00040, 16'd00040, 16'd00000, 16'd00040, 16'd00080, 16'd000C1, 16'd00101, 16'd000C0, 16'd00000, 16'd00000, 16'd00040, 16'd06247, 16'd13594, 16'd1F921, 16'd27B2A, 16'd25AA7, 16'd1B7DD, 16'd0E44F, 16'd03143, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd03000, 16'd03000, 16'd03000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00080, 16'd00080, 16'd00080, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00080, 16'd000C1, 16'd00101, 16'd000C0, 16'd00000, 16'd00000, 16'd00040, 16'd06247, 16'd13594, 16'd20922, 16'd27B2A, 16'd25AA8, 16'd1B7DD, 16'd0E44F, 16'd03143, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00080, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00080, 16'd000C1, 16'd000C1, 16'd00080, 16'd00000, 16'd00000, 16'd00040, 16'd07247, 16'd135D5, 16'd20962, 16'd28B6B, 16'd26AE9, 16'd1C81E, 16'd0E44F, 16'd03143, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00080, 16'd00081, 16'd000C1, 16'd000C1, 16'd00080, 16'd00000, 16'd00000, 16'd00040, 16'd07247, 16'd145D5, 16'd229A4, 16'd2ABED, 16'd28B2A, 16'd1D85F, 16'd0F490, 16'd03143, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd01040, 16'd01040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00080, 16'd00080, 16'd00081, 16'd000C1, 16'd000C1, 16'd000C1, 16'd00080, 16'd00000, 16'd00000, 16'd00000, 16'd07247, 16'd15616, 16'd239E5, 16'd2CC2E, 16'd29BAC, 16'd1E8A0, 16'd0F490, 16'd03143, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd01040, 16'd01040, 16'd01040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00081, 16'd01081, 16'd010C1, 16'd000C1, 16'd000C1, 16'd000C0, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd07247, 16'd16657, 16'd24A26, 16'd2DCAF, 16'd2BBED, 16'd1F8E1, 16'd104D1, 16'd03143, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01040, 16'd01040, 16'd01040, 16'd01040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd01081, 16'd010C1, 16'd010C1, 16'd000C1, 16'd00080, 16'd00080, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd07248, 16'd16657, 16'd25A67, 16'd2ECB0, 16'd2CC2E, 16'd208E1, 16'd104D1, 16'd03143, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01040, 16'd01040, 16'd01040, 16'd01040, 16'd01040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd01081, 16'd01081, 16'd01081, 16'd00080, 16'd00080, 16'd00080, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd08288, 16'd16657, 16'd25A67, 16'd2ECB0, 16'd2CC2E, 16'd208E1, 16'd104D1, 16'd03143, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01040, 16'd01040, 16'd01040, 16'd01040, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd01040, 16'd01040, 16'd01081, 16'd00080, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd08288, 16'd17698, 16'd26A67, 16'd2FCB0, 16'd2CC2E, 16'd208E2, 16'd104D1, 16'd03143, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01040, 16'd01040, 16'd01040, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd082C9, 16'd17698, 16'd26A67, 16'd2ECB0, 16'd2CBEE, 16'd208E1, 16'd10491, 16'd03143, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd02040, 16'd02040, 16'd02040, 16'd02040, 16'd02000, 16'd02040, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00080, 16'd082C9, 16'd16657, 16'd25A26, 16'd2DC2F, 16'd2BBAC, 16'd1F8A0, 16'd10490, 16'd03143, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd02000, 16'd02040, 16'd02040, 16'd02040, 16'd02040, 16'd02040, 16'd02040, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00080, 16'd07288, 16'd15616, 16'd22963, 16'd2AB6B, 16'd28AE9, 16'd1D7DE, 16'd0F44F, 16'd03103, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd02000, 16'd02040, 16'd02040, 16'd02040, 16'd02040, 16'd02040, 16'd02040, 16'd02040, 16'd02040, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00080, 16'd06247, 16'd12553, 16'd1D81E, 16'd249E5, 16'd22963, 16'd196DA, 16'd0D3CD, 16'd02102, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd02041, 16'd02041, 16'd03041, 16'd02041, 16'd02040, 16'd02040, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd01040, 16'd01041, 16'd01041, 16'd01041, 16'd00040, 16'd00000, 16'd00040, 16'd051C5, 16'd0D40E, 16'd16657, 16'd1C79D, 16'd1A75B, 16'd13554, 16'd0A2CA, 16'd020C2, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01041, 16'd03082, 16'd040C2, 16'd040C2, 16'd03082, 16'd03041, 16'd02040, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd01040, 16'd02041, 16'd02081, 16'd020C2, 16'd02081, 16'd01041, 16'd00000, 16'd00040, 16'd03103, 16'd08289, 16'd0E44F, 16'd12513, 16'd114D2, 16'd0C3CD, 16'd06206, 16'd010C1, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd02041, 16'd030C2, 16'd05103, 16'd05103, 16'd040C2, 16'd03081, 16'd02040, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01040, 16'd02081, 16'd030C2, 16'd03102, 16'd030C2, 16'd01081, 16'd00000, 16'd00000, 16'd01081, 16'd04144, 16'd07248, 16'd092CA, 16'd082C9, 16'd06207, 16'd03143, 16'd00080, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd02081, 16'd040C3, 16'd05104, 16'd06144, 16'd04103, 16'd03081, 16'd01040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01040, 16'd02080, 16'd030C1, 16'd03102, 16'd04103, 16'd03102, 16'd02081, 16'd01040, 16'd00000, 16'd00040, 16'd00081, 16'd010C2, 16'd02103, 16'd02103, 16'd010C2, 16'd00081, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd02081, 16'd040C2, 16'd05103, 16'd05104, 16'd040C3, 16'd03081, 16'd01040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01040, 16'd02080, 16'd020C1, 16'd030C2, 16'd03103, 16'd03102, 16'd020C1, 16'd01041, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01041, 16'd03082, 16'd040C3, 16'd040C3, 16'd030C2, 16'd02041, 16'd01040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01040, 16'd01040, 16'd02081, 16'd020C2, 16'd030C2, 16'd020C2, 16'd020C1, 16'd01081, 16'd01041, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01040, 16'd02041, 16'd02081, 16'd03082, 16'd02081, 16'd01040, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd01040, 16'd01040, 16'd01081, 16'd02081, 16'd02081, 16'd020C1, 16'd020C2, 16'd020C1, 16'd01081, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01040, 16'd01040, 16'd01040, 16'd01040, 16'd00040, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd01040, 16'd01081, 16'd010C1, 16'd020C2, 16'd02102, 16'd020C2, 16'd01081, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd01081, 16'd02102, 16'd03103, 16'd02102, 16'd020C2, 16'd01041, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00080, 16'd00080, 16'd00080, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd01081, 16'd020C2, 16'd02102, 16'd02102, 16'd020C1, 16'd01040, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd01081, 16'd010C1, 16'd020C2, 16'd020C2, 16'd01081, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00040, 16'd00040, 16'd01081, 16'd01081, 16'd01081, 16'd01040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00080, 16'd000C1, 16'd000C0, 16'd000C0, 16'd00080, 16'd00040, 16'd00040, 16'd00040, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd010C2, 16'd02184, 16'd03205, 16'd03246, 16'd03246, 16'd03205, 16'd031C4, 16'd031C3, 16'd031C3, 16'd031C4, 16'd031C4, 16'd031C4, 16'd02183, 16'd01142, 16'd00101, 16'd000C0, 16'd000C0, 16'd00080, 16'd00080, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01081, 16'd041C5, 16'd0730A, 16'd0A44D, 16'd0B4CF, 16'd0B4CF, 16'd0B44E, 16'd0A40C, 16'd0A40C, 16'd0A40C, 16'd0A44D, 16'd0A44D, 16'd0940C, 16'd0734A, 16'd04287, 16'd011C4, 16'd00141, 16'd000C0, 16'd00080, 16'd00080, 16'd00040, 16'd00040, 16'd00040, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00081, 16'd00081, 16'd00041, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd020C2, 16'd072C9, 16'd0D4D0, 16'd13697, 16'd1579A, 16'd1579A, 16'd14759, 16'd13717, 16'd126D6, 16'd136D7, 16'd13717, 16'd13717, 16'd12696, 16'd0E591, 16'd0840C, 16'd032C7, 16'd001C3, 16'd00101, 16'd000C0, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd000C1, 16'd000C1, 16'd000C1, 16'd000C1, 16'd010C1, 16'd00081, 16'd00081, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd02103, 16'd0A38C, 16'd14697, 16'd1B920, 16'd1FA64, 16'd1FAA5, 16'd1DA23, 16'd1B9E1, 16'd1B9A0, 16'd1B9A1, 16'd1C9E2, 16'd1C9A2, 16'd1A91F, 16'd14799, 16'd0C591, 16'd0438A, 16'd00204, 16'd00141, 16'd000C0, 16'd000C0, 16'd00080, 16'd00080, 16'd00080, 16'd000C1, 16'd00101, 16'd00101, 16'd00102, 16'd01102, 16'd01102, 16'd010C2, 16'd00081, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd03144, 16'd0D48F, 16'd1981C, 16'd23B28, 16'd27CAD, 16'd27CEE, 16'd25C6C, 16'd22BE9, 16'd21BA8, 16'd22BE9, 16'd23C2A, 16'd23BEA, 16'd20B27, 16'd1991F, 16'd0F696, 16'd0640C, 16'd00245, 16'd00141, 16'd00100, 16'd000C0, 16'd00080, 16'd00080, 16'd000C0, 16'd00101, 16'd00102, 16'd00142, 16'd00142, 16'd01143, 16'd01143, 16'd01102, 16'd010C2, 16'd00041, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd04184, 16'd0F511, 16'd1C920, 16'd27C6D, 16'd2CE33, 16'd2CE73, 16'd29DF1, 16'd26D2E, 16'd24CED, 16'd26D2E, 16'd27D6F, 16'd27D6F, 16'd24C6C, 16'd1CA23, 16'd11758, 16'd0644C, 16'd00245, 16'd00141, 16'd000C0, 16'd000C0, 16'd000C0, 16'd000C0, 16'd000C0, 16'd00101, 16'd00142, 16'd00142, 16'd00142, 16'd01142, 16'd01102, 16'd01102, 16'd010C2, 16'd00081, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd041C5, 16'd10553, 16'd1E9E3, 16'd2AD70, 16'd2FF37, 16'd2FF77, 16'd2BEB3, 16'd27DB0, 16'd25D6E, 16'd27DB0, 16'd29E31, 16'd29E32, 16'd26D2E, 16'd1EAA5, 16'd12758, 16'd0744C, 16'd00204, 16'd00101, 16'd000C0, 16'd000C0, 16'd000C0, 16'd000C0, 16'd000C0, 16'd00101, 16'd00141, 16'd00141, 16'd00102, 16'd00102, 16'd01102, 16'd010C2, 16'd010C2, 16'd01081, 16'd01081, 16'd01041, 16'd01041, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd041C5, 16'd115D4, 16'd20A25, 16'd2CE33, 16'd31FB9, 16'd30FB8, 16'd2BEF4, 16'd27DF0, 16'd25D6E, 16'd26DF0, 16'd29E72, 16'd2AE73, 16'd27D6F, 16'd1EAE6, 16'd13758, 16'd0740B, 16'd001C2, 16'd000C1, 16'd00080, 16'd000C0, 16'd000C0, 16'd000C0, 16'd00100, 16'd00100, 16'd00101, 16'd00101, 16'd000C1, 16'd000C1, 16'd000C1, 16'd00081, 16'd01081, 16'd010C2, 16'd020C2, 16'd02082, 16'd01081, 16'd01040, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd041C5, 16'd125D4, 16'd21AA6, 16'd2DE74, 16'd32FFA, 16'd30FF9, 16'd2BEF4, 16'd26DAF, 16'd24D6D, 16'd25DAF, 16'd28E72, 16'd2AEB3, 16'd27DB0, 16'd1FAE6, 16'd13758, 16'd073CA, 16'd00141, 16'd00080, 16'd00080, 16'd000C0, 16'd00100, 16'd00100, 16'd00100, 16'd00100, 16'd00100, 16'd000C0, 16'd000C0, 16'd00080, 16'd00040, 16'd00080, 16'd01081, 16'd020C2, 16'd02103, 16'd03103, 16'd02082, 16'd01041, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd041C5, 16'd12614, 16'd21AA6, 16'd2DEB5, 16'd32FFB, 16'd30FF9, 16'd2BEF4, 16'd25DAF, 16'd23D2D, 16'd25DAF, 16'd28E72, 16'd29EB3, 16'd27DB0, 16'd1EAE5, 16'd13717, 16'd07389, 16'd00100, 16'd00040, 16'd00040, 16'd000C0, 16'd00100, 16'd00100, 16'd00100, 16'd00100, 16'd000C0, 16'd000C0, 16'd00080, 16'd00040, 16'd00040, 16'd00040, 16'd01081, 16'd02103, 16'd03144, 16'd03103, 16'd030C3, 16'd02081, 16'd01000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd041C5, 16'd12614, 16'd21AA6, 16'd2DEB5, 16'd32FFB, 16'd30FF9, 16'd2AEF4, 16'd25DAF, 16'd23D2D, 16'd24DAF, 16'd28E72, 16'd29EB4, 16'd27DB0, 16'd1EAE5, 16'd13717, 16'd07349, 16'd00100, 16'd00040, 16'd00040, 16'd000C0, 16'd00100, 16'd00100, 16'd00100, 16'd000C0, 16'd000C0, 16'd000C0, 16'd00080, 16'd00040, 16'd00040, 16'd00080, 16'd010C2, 16'd02103, 16'd03144, 16'd03103, 16'd030C3, 16'd02081, 16'd01000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd041C5, 16'd115D4, 16'd20AA6, 16'd2CE74, 16'd31FFA, 16'd30FF9, 16'd2BF35, 16'd25DF0, 16'd23DAE, 16'd25DF0, 16'd28EB3, 16'd2AEF4, 16'd27DB0, 16'd1EAE5, 16'd13717, 16'd07389, 16'd00100, 16'd00040, 16'd00040, 16'd000C0, 16'd00100, 16'd00100, 16'd00100, 16'd000C0, 16'd000C0, 16'd000C0, 16'd00080, 16'd01081, 16'd010C1, 16'd010C2, 16'd020C2, 16'd02103, 16'd03103, 16'd030C3, 16'd02082, 16'd01041, 16'd01000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd01000, 16'd01000, 16'd01000, 16'd01000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd041C5, 16'd115D3, 16'd1FA64, 16'd2BE33, 16'd30FF9, 16'd2FFF9, 16'd2BF35, 16'd26E31, 16'd24DEF, 16'd26E71, 16'd28EB3, 16'd29EF4, 16'd27DB0, 16'd1EAE5, 16'd12757, 16'd07389, 16'd00140, 16'd00040, 16'd00040, 16'd000C0, 16'd00100, 16'd00100, 16'd000C0, 16'd000C0, 16'd00080, 16'd000C0, 16'd010C1, 16'd02102, 16'd03143, 16'd03143, 16'd03103, 16'd020C3, 16'd020C2, 16'd02082, 16'd01081, 16'd01040, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd01000, 16'd01000, 16'd01000, 16'd01000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd041C5, 16'd10592, 16'd1D9E3, 16'd28DB0, 16'd2DF77, 16'd2DFB7, 16'd2AF34, 16'd26E71, 16'd25DF0, 16'd26E71, 16'd28EB3, 16'd29EB3, 16'd25D6F, 16'd1DAE4, 16'd12717, 16'd073C9, 16'd00180, 16'd00080, 16'd00080, 16'd000C0, 16'd00100, 16'd000C0, 16'd000C0, 16'd00080, 16'd00080, 16'd000C0, 16'd02102, 16'd03184, 16'd041C5, 16'd04185, 16'd03144, 16'd020C3, 16'd01081, 16'd01041, 16'd00041, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd01000, 16'd01000, 16'd01000, 16'd01000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd04184, 16'd0E511, 16'd1B920, 16'd25CAC, 16'd2AE73, 16'd2AEB4, 16'd28E72, 16'd25DEF, 16'd24DAE, 16'd25DF0, 16'd26E31, 16'd26DF0, 16'd23CED, 16'd1BA63, 16'd11716, 16'd063C9, 16'd00181, 16'd00080, 16'd00080, 16'd000C0, 16'd00100, 16'd000C0, 16'd000C0, 16'd00080, 16'd00080, 16'd010C1, 16'd02143, 16'd04185, 16'd05206, 16'd051C6, 16'd03144, 16'd020C2, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd03184, 16'd0C48F, 16'd1781C, 16'd20B27, 16'd25CED, 16'd25D2E, 16'd23CEC, 16'd21CAA, 16'd20C6A, 16'd21CAB, 16'd22CEC, 16'd22CAC, 16'd1FBA8, 16'd1895F, 16'd0F653, 16'd05388, 16'd00181, 16'd000C0, 16'd00080, 16'd000C0, 16'd00100, 16'd000C0, 16'd00080, 16'd00080, 16'd00080, 16'd010C1, 16'd02103, 16'd04185, 16'd05206, 16'd051C6, 16'd03144, 16'd01082, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd02143, 16'd0A3CC, 16'd12696, 16'd1991F, 16'd1DA63, 16'd1DAA4, 16'd1CAA3, 16'd1AA62, 16'd1AA21, 16'd1AAA3, 16'd1BAA4, 16'd1BAA4, 16'd199E1, 16'd1381A, 16'd0B590, 16'd04307, 16'd00180, 16'd000C0, 16'd00080, 16'd000C0, 16'd000C0, 16'd000C0, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd02102, 16'd03144, 16'd04185, 16'd04185, 16'd03103, 16'd01081, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01102, 16'd062C8, 16'd0C4CF, 16'd11655, 16'd13758, 16'd14799, 16'd13798, 16'd12757, 16'd11757, 16'd127D8, 16'd1281A, 16'd1281A, 16'd11799, 16'd0D653, 16'd0844C, 16'd03285, 16'd00140, 16'd00080, 16'd00080, 16'd000C0, 16'd000C0, 16'd00080, 16'd00080, 16'd00040, 16'd00040, 16'd00080, 16'd010C1, 16'd02103, 16'd03144, 16'd03103, 16'd020C2, 16'd00041, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01081, 16'd031C4, 16'd062C8, 16'd093CB, 16'd0A48D, 16'd0A48D, 16'd0A48D, 16'd0948C, 16'd0948C, 16'd0950E, 16'd0A550, 16'd0A591, 16'd09590, 16'd0748C, 16'd04348, 16'd011C3, 16'd00100, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00040, 16'd00040, 16'd00040, 16'd00081, 16'd01081, 16'd010C2, 16'd01082, 16'd01041, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00080, 16'd010C1, 16'd02142, 16'd021C3, 16'd03203, 16'd03203, 16'd03203, 16'd02203, 16'd02243, 16'd02285, 16'd02307, 16'd02388, 16'd02388, 16'd02307, 16'd01244, 16'd00141, 16'd000C0, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd000C0, 16'd00140, 16'd001C2, 16'd00203, 16'd00244, 16'd00203, 16'd00182, 16'd00101, 16'd000C0, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00080, 16'd00100, 16'd00141, 16'd00181, 16'd00181, 16'd00141, 16'd00100, 16'd000C0, 16'd000C0, 16'd000C0, 16'd000C0, 16'd000C0, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00080, 16'd000C0, 16'd00100, 16'd00100, 16'd00101, 16'd00101, 16'd00101, 16'd00101, 16'd00101, 16'd00101, 16'd000C1, 16'd000C1, 16'd010C1, 16'd010C1, 16'd010C1, 16'd01081, 16'd00080, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01041, 16'd01041, 16'd01041, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00080, 16'd00080, 16'd000C0, 16'd000C0, 16'd00100, 16'd00101, 16'd00101, 16'd00101, 16'd00101, 16'd00102, 16'd01102, 16'd01102, 16'd01102, 16'd01101, 16'd010C1, 16'd010C1, 16'd01081, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01041, 16'd02081, 16'd02081, 16'd02041, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd00000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd000C0, 16'd000C0, 16'd000C0, 16'd00101, 16'd00101, 16'd00102, 16'd00142, 16'd00142, 16'd01142, 16'd01102, 16'd01102, 16'd01102, 16'd01102, 16'd010C1, 16'd01081, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd01040, 16'd02081, 16'd02082, 16'd02082, 16'd02081, 16'd01041, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd000C1, 16'd00101, 16'd00102, 16'd00142, 16'd00142, 16'd01142, 16'd01102, 16'd01102, 16'd01102, 16'd01102, 16'd010C1, 16'd01081, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd01040, 16'd02081, 16'd03082, 16'd03082, 16'd02081, 16'd01041, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00040, 16'd00040, 16'd00040, 16'd00080, 16'd00080, 16'd000C1, 16'd00101, 16'd00102, 16'd00102, 16'd01102, 16'd01102, 16'd010C2, 16'd010C2, 16'd010C1, 16'd01081, 16'd01081, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd02041, 16'd02082, 16'd02082, 16'd02041, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00080, 16'd00080, 16'd00080, 16'd000C0, 16'd00080, 16'd00080, 16'd00080, 16'd00080, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00080, 16'd00080, 16'd000C1, 16'd000C1, 16'd000C1, 16'd000C1, 16'd00081, 16'd01081, 16'd01081, 16'd01081, 16'd01081, 16'd01041, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01041, 16'd02041, 16'd02041, 16'd01041, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00080, 16'd00081, 16'd000C1, 16'd000C0, 16'd000C0, 16'd00080, 16'd00080, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00080, 16'd00080, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01040, 16'd01040, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00080, 16'd00080, 16'd00080, 16'd00080,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00081, 16'd000C1, 16'd000C1, 16'd000C1, 16'd00080, 16'd00080, 16'd00080, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00080, 16'd00080, 16'd00080, 16'd00080,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00081, 16'd000C1, 16'd000C1, 16'd000C1, 16'd00080, 16'd00080, 16'd00080, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00080, 16'd00080, 16'd00080, 16'd00080,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00081, 16'd00081, 16'd00080, 16'd00080, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00080, 16'd00080, 16'd00080, 16'd00080,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00080, 16'd00080, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02041, 16'd02001, 16'd01000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00080, 16'd00080, 16'd00080, 16'd00080,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02040, 16'd02041, 16'd02041, 16'd02041, 16'd02041, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00080, 16'd00080, 16'd00080, 16'd00080,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02040, 16'd02041, 16'd03041, 16'd03082, 16'd03042, 16'd02041, 16'd02000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02040, 16'd02041, 16'd03041, 16'd03082, 16'd03042, 16'd02041, 16'd02000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02040, 16'd02040, 16'd02040, 16'd02040, 16'd02000, 16'd02000, 16'd02000, 16'd02040, 16'd03041, 16'd03041, 16'd03041, 16'd02041, 16'd01000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02040, 16'd03041, 16'd03081, 16'd03041, 16'd02040, 16'd02040, 16'd01000, 16'd01000, 16'd02040, 16'd02041, 16'd02041, 16'd02041, 16'd02000, 16'd01000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02040, 16'd02041, 16'd03081, 16'd03081, 16'd03081, 16'd02041, 16'd02040, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02040, 16'd03041, 16'd04082, 16'd040C2, 16'd03082, 16'd02081, 16'd01040, 16'd01000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02040, 16'd03081, 16'd040C2, 16'd040C2, 16'd03082, 16'd02081, 16'd01040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02040, 16'd02081, 16'd030C2, 16'd040C2, 16'd03082, 16'd02081, 16'd01040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01040, 16'd02081, 16'd030C2, 16'd030C2, 16'd03082, 16'd02081, 16'd01040, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01040, 16'd02081, 16'd02081, 16'd030C2, 16'd02081, 16'd01041, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01041, 16'd01041, 16'd01040, 16'd01040, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd01041, 16'd02081, 16'd02081, 16'd02081, 16'd01041, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01040, 16'd01041, 16'd01041, 16'd01041, 16'd01041, 16'd01040, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd01040, 16'd01081, 16'd02081, 16'd01081, 16'd01040, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd01041, 16'd02081, 16'd02081, 16'd02041, 16'd01041, 16'd01040, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd01040, 16'd01080, 16'd01081, 16'd01080, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd01041, 16'd02081, 16'd02081, 16'd02041, 16'd01041, 16'd01040, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00080, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd01040, 16'd01040, 16'd01040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd01041, 16'd02081, 16'd02081, 16'd01041, 16'd01040, 16'd01000, 16'd01000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00080, 16'd01081, 16'd01081, 16'd00081, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd01081, 16'd02081, 16'd02081, 16'd01041, 16'd01040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd01081, 16'd010C1, 16'd010C1, 16'd010C1, 16'd00080, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd01081, 16'd01081, 16'd01081, 16'd01041, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00080, 16'd010C1, 16'd010C1, 16'd01101, 16'd010C1, 16'd00080, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd01081, 16'd01081, 16'd01081, 16'd01041, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00080, 16'd010C1, 16'd01102, 16'd01102, 16'd010C1, 16'd00080, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd01081, 16'd01081, 16'd01081, 16'd01041, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000,
        16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd00080, 16'd010C1, 16'd01102, 16'd01102, 16'd010C1, 16'd00080, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00040, 16'd00040, 16'd00040, 16'd00040, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00040, 16'd01081, 16'd01081, 16'd01081, 16'd01041, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd00000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd01000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd02000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd03000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000, 16'd04000,
    };
    reg [0:15] img_out [21384:0];

    always @(*) begin
        if(step == 0) img_out <= step0;
        else img_out <= img_out;
    end

    integer i;
    always @(*) begin
        for(i = 0; i < 132; i = i + 1) begin
            ram_data[i] <= img_out[ram_addr * 132 + i];
        end
    end
    
endmodule