module idle_mem (
    input [3:0] step,
    input [7:0] ram_addr_x,
    input [7:0] ram_addr_y,
    output reg[15:0] ram_data
);

    parameter [15:0] step0 [0:131] = {
        16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0020, 16'h0040, 16'h0060, 16'h0081, 16'h0081, 16'h0060, 16'h0040, 16'h0020, 16'h0020, 16'h0000, 16'h0000, 16'h0020, 16'h0020, 16'h0020, 16'h0020, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0020, 16'h0040, 16'h0040, 16'h0040, 16'h0020, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0800, 16'h0800, 16'h0800, 16'h0800, 16'h0800, 16'h0800, 16'h0800, 16'h0800, 16'h0800, 16'h0800, 16'h0800, 16'h0800, 16'h0800, 16'h0800, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000
    };

    always @(*) begin
        if(step == 0) ram_data = step0[ram_addr_y*132 + ram_addr_x];
    end
    
endmodule