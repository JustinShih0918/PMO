module idle_mem (
    input [3:0] step,
    input [7:0] ram_addr_x,
    input [7:0] ram_addr_y,
    output [15:0] ram_data
);

    parameter [0:15] step0 [21384:0] = {
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0040, 16'd0060, 16'd0081, 16'd0081, 16'd0060, 16'd0040, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0040, 16'd0060, 16'd0081, 16'd0081, 16'd0060, 16'd0040, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0040, 16'd0060, 16'd0060, 16'd0080, 16'd0060, 16'd0040, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0040, 16'd0040, 16'd0060, 16'd0060, 16'd0060, 16'd0040, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0040, 16'd0840, 16'd0840, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0840, 16'd0840, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0840, 16'd0840, 16'd0820, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0040, 16'd0840, 16'd0040, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0840, 16'd0840, 16'd0820, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0840, 16'd0840, 16'd0840, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0840, 16'd0840, 16'd0861, 16'd0840, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0840, 16'd0861, 16'd0861, 16'd0841, 16'd0840, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0820, 16'd0840, 16'd0861, 16'd1061, 16'd0841, 16'd0840, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0820, 16'd0840, 16'd1061, 16'd1061, 16'd0841, 16'd0840, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0820, 16'd0820, 16'd1041, 16'd1061, 16'd0841, 16'd0840, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0820, 16'd0820, 16'd0840, 16'd0840, 16'd0840, 16'd0820, 16'd0820, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0820, 16'd0820, 16'd0840, 16'd0820, 16'd0820, 16'd0820, 16'd0000, 16'd0000, 16'd0820, 16'd0820, 16'd0820, 16'd0820, 16'd0800, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0820, 16'd0820, 16'd0820, 16'd0820, 16'd0800, 16'd0800, 16'd0800, 16'd0820, 16'd0820, 16'd0820, 16'd0820, 16'd0820, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0820, 16'd0820, 16'd0820, 16'd0841, 16'd0821, 16'd0820, 16'd0800, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0820, 16'd0820, 16'd0820, 16'd0841, 16'd0821, 16'd0820, 16'd0800, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0820, 16'd0820, 16'd0820, 16'd0820, 16'd0820, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0040,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0820, 16'd0800, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0040,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0040,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0040, 16'd0060, 16'd0060, 16'd0060, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0040,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0040, 16'd0060, 16'd0060, 16'd0060, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0040,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0040, 16'd0040, 16'd0060, 16'd0060, 16'd0060, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0040,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0060, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0060, 16'd0060, 16'd0060, 16'd0060, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0820, 16'd0820, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0060, 16'd0080, 16'd0081, 16'd0081, 16'd0081, 16'd0081, 16'd0061, 16'd0061, 16'd0060, 16'd0040, 16'd0040, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0820, 16'd0841, 16'd0841, 16'd0820, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0060, 16'd0080, 16'd0081, 16'd00A1, 16'd00A1, 16'd00A1, 16'd0081, 16'd0081, 16'd0081, 16'd0081, 16'd0060, 16'd0040, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0840, 16'd0841, 16'd0841, 16'd0840, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0060, 16'd0060, 16'd0060, 16'd0080, 16'd0080, 16'd0081, 16'd00A1, 16'd00A1, 16'd00A1, 16'd0081, 16'd0081, 16'd0081, 16'd0081, 16'd0060, 16'd0040, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0840, 16'd0841, 16'd0841, 16'd0840, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0060, 16'd0060, 16'd0080, 16'd0080, 16'd0080, 16'd0080, 16'd0080, 16'd0081, 16'd0081, 16'd0081, 16'd0081, 16'd0080, 16'd0060, 16'd0060, 16'd0040, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0840, 16'd0840, 16'd0820, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0040, 16'd0060, 16'd0080, 16'd0080, 16'd0080, 16'd0080, 16'd0080, 16'd0080, 16'd0080, 16'd0080, 16'd0060, 16'd0060, 16'd0060, 16'd0060, 16'd0060, 16'd0040, 16'd0040, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0040, 16'd0080, 16'd00A0, 16'd00C0, 16'd00C0, 16'd00A0, 16'd0080, 16'd0060, 16'd0060, 16'd0060, 16'd0060, 16'd0060, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0060, 16'd00A0, 16'd00E1, 16'd0101, 16'd0122, 16'd0101, 16'd00C1, 16'd0080, 16'd0060, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0040, 16'd0060, 16'd08A1, 16'd08E1, 16'd0901, 16'd0901, 16'd0901, 16'd0901, 16'd0921, 16'd0942, 16'd0983, 16'd09C4, 16'd09C4, 16'd0983, 16'd0122, 16'd00A0, 16'd0060, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0040, 16'd08E2, 16'd1964, 16'd21E5, 16'd2A46, 16'd2A46, 16'd2A46, 16'd2246, 16'd2246, 16'd2287, 16'd2AA8, 16'd2AC8, 16'd22C8, 16'd1A46, 16'd11A4, 16'd00E1, 16'd0080, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0061, 16'd0041, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0081, 16'd1964, 16'd3267, 16'd432A, 16'd4BAC, 16'd53CC, 16'd4BCC, 16'd4BAB, 16'd43AB, 16'd4BEC, 16'd4C0D, 16'd4C0D, 16'd43CC, 16'd3329, 16'd2226, 16'd0942, 16'd00A0, 16'd0040, 16'd0040, 16'd0060, 16'd0060, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0040, 16'd0060, 16'd0881, 16'd08A2, 16'd0881, 16'd0861, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd08A1, 16'd29E6, 16'd4B4B, 16'd648F, 16'd7531, 16'd7552, 16'd7551, 16'd6D31, 16'd6D10, 16'd6D51, 16'd6D52, 16'd6D52, 16'd64F0, 16'd4C0D, 16'd2AC8, 16'd1183, 16'd00C0, 16'd0060, 16'd0040, 16'd0060, 16'd0060, 16'd0060, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0881, 16'd08A2, 16'd10C2, 16'd10C2, 16'd0881, 16'd0040, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd08C2, 16'd3247, 16'd5C0E, 16'd8593, 16'd9676, 16'd9697, 16'd8E76, 16'd8655, 16'd8635, 16'd8655, 16'd8E76, 16'd8E56, 16'd7DD4, 16'd64AF, 16'd3B29, 16'd11C4, 16'd00C0, 16'd0060, 16'd0040, 16'd0060, 16'd0080, 16'd0060, 16'd0040, 16'd0040, 16'd0040, 16'd0060, 16'd0881, 16'd10C2, 16'd1103, 16'd10E3, 16'd08A2, 16'd0041, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd10C2, 16'd3A88, 16'd6C90, 16'd9656, 16'dAF39, 16'dAF5A, 16'dA739, 16'd96F7, 16'd96D7, 16'd96F8, 16'd9F18, 16'd9EF8, 16'd8E76, 16'd6D31, 16'd438B, 16'd19E4, 16'd00C0, 16'd0040, 16'd0040, 16'd0060, 16'd0080, 16'd0060, 16'd0060, 16'd0040, 16'd0040, 16'd0060, 16'd08A1, 16'd10C2, 16'd1103, 16'd10E3, 16'd08A2, 16'd0861, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd10E2, 16'd42C9, 16'd74F1, 16'dA6D8, 16'dB7BB, 16'dB7DB, 16'dAF9A, 16'd9F38, 16'd96F8, 16'd9F38, 16'dA759, 16'dA759, 16'd96B7, 16'd7572, 16'd4B8B, 16'd19E4, 16'd00C0, 16'd0040, 16'd0040, 16'd0060, 16'd0080, 16'd0060, 16'd0060, 16'd0040, 16'd0040, 16'd0060, 16'd0881, 16'd08C2, 16'd10E2, 16'd10C2, 16'd08A2, 16'd0861, 16'd0040, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd10E2, 16'd42E9, 16'd7D32, 16'dAF19, 16'dC7FC, 16'dBFFC, 16'dAF9A, 16'd9F18, 16'd96F7, 16'd9F38, 16'dA759, 16'dA77A, 16'd9ED8, 16'd7D72, 16'd4BAB, 16'd19C4, 16'd00A0, 16'd0020, 16'd0020, 16'd0060, 16'd0080, 16'd0080, 16'd0060, 16'd0060, 16'd0040, 16'd0060, 16'd0060, 16'd0881, 16'd08A1, 16'd08A1, 16'd0881, 16'd0861, 16'd0861, 16'd0841, 16'd0040, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd10E2, 16'd42EA, 16'd8553, 16'dB73A, 16'dC7FD, 16'dC7FC, 16'dAF9A, 16'd96F8, 16'd8ED7, 16'd96F8, 16'dA759, 16'dAF7A, 16'd9ED8, 16'd7D72, 16'd4B8B, 16'd19C4, 16'd0080, 16'd0020, 16'd0020, 16'd0060, 16'd0080, 16'd0080, 16'd0080, 16'd0060, 16'd0060, 16'd0060, 16'd0040, 16'd0040, 16'd0060, 16'd0061, 16'd0861, 16'd0881, 16'd0881, 16'd0861, 16'd0841, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd10E2, 16'd4B0A, 16'd8553, 16'dB75A, 16'dCFFD, 16'dC7FC, 16'dAF7A, 16'd96D7, 16'd8E96, 16'd96D7, 16'dA739, 16'dA75A, 16'd9ED8, 16'd7D72, 16'd4B8B, 16'd19A4, 16'd0080, 16'd0020, 16'd0020, 16'd0060, 16'd0080, 16'd0080, 16'd0080, 16'd0060, 16'd0060, 16'd0060, 16'd0040, 16'd0020, 16'd0020, 16'd0040, 16'd0061, 16'd0881, 16'd08A2, 16'd0881, 16'd0861, 16'd0840, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd10E2, 16'd4B0A, 16'd8553, 16'dB75A, 16'dCFFD, 16'dC7FC, 16'dAF7A, 16'd96D7, 16'd8E96, 16'd96D7, 16'dA739, 16'dA759, 16'd9ED8, 16'd7D72, 16'd4B8B, 16'd19C4, 16'd0080, 16'd0020, 16'd0020, 16'd0060, 16'd0080, 16'd0080, 16'd0080, 16'd0080, 16'd0060, 16'd0060, 16'd0040, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0881, 16'd08A2, 16'd0881, 16'd0861, 16'd0840, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd10E2, 16'd4AEA, 16'd8553, 16'dB73A, 16'dCFFD, 16'dC7FC, 16'dAF7A, 16'd9ED7, 16'd96B6, 16'd96D7, 16'dA739, 16'dAF59, 16'd9ED8, 16'd7D73, 16'd4BAC, 16'd19E5, 16'd00A0, 16'd0040, 16'd0040, 16'd0060, 16'd0080, 16'd0080, 16'd0080, 16'd0080, 16'd0080, 16'd0060, 16'd0060, 16'd0040, 16'd0020, 16'd0040, 16'd0040, 16'd0861, 16'd0881, 16'd0881, 16'd0841, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd10E2, 16'd42EA, 16'd8512, 16'dB719, 16'dC7DC, 16'dC7DC, 16'dAF7A, 16'd9EF8, 16'd96B7, 16'd9EF8, 16'dA739, 16'dAF39, 16'd9EB7, 16'd7D73, 16'd4BAC, 16'd1A05, 16'd00E1, 16'd0060, 16'd0040, 16'd0060, 16'd0060, 16'd0060, 16'd0080, 16'd0080, 16'd0080, 16'd0080, 16'd0060, 16'd0060, 16'd0060, 16'd0040, 16'd0040, 16'd0061, 16'd0861, 16'd0841, 16'd0040, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd10E2, 16'd42A9, 16'd7CF1, 16'dAEB8, 16'dBF9B, 16'dBFBB, 16'dAF59, 16'd9ED8, 16'd96B7, 16'd9ED8, 16'dA718, 16'dA719, 16'd9E97, 16'd7D52, 16'd4BAC, 16'd1A26, 16'd0102, 16'd0080, 16'd0060, 16'd0060, 16'd0060, 16'd0060, 16'd0060, 16'd0080, 16'd00A0, 16'd00A0, 16'd0081, 16'd0081, 16'd0081, 16'd0061, 16'd0061, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd10C2, 16'd3A88, 16'd7490, 16'd9E36, 16'dB719, 16'dB739, 16'dA6F8, 16'd9E97, 16'd9676, 16'd9E97, 16'd9EB7, 16'd9EB7, 16'd9636, 16'd7511, 16'd43AC, 16'd1A26, 16'd0122, 16'd00A0, 16'd0060, 16'd0060, 16'd0060, 16'd0060, 16'd0060, 16'd0080, 16'd00A1, 16'd00A1, 16'd00A1, 16'd00A1, 16'd0081, 16'd0081, 16'd0061, 16'd0040, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd08A2, 16'd3247, 16'd640E, 16'd8D94, 16'd9E56, 16'd9E77, 16'd9636, 16'd8DF4, 16'd85D4, 16'd8DF4, 16'd8E15, 16'd8DF5, 16'd8593, 16'd648F, 16'd3B4B, 16'd1A06, 16'd0122, 16'd00A0, 16'd0080, 16'd0060, 16'd0040, 16'd0040, 16'd0060, 16'd0080, 16'd0081, 16'd00A1, 16'd00A1, 16'd00A1, 16'd00A1, 16'd0081, 16'd0061, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0881, 16'd29C6, 16'd534B, 16'd6C90, 16'd7D32, 16'd7D52, 16'd7511, 16'd6CF0, 16'd6CD0, 16'd6CD0, 16'd74F1, 16'd74D1, 16'd6C8F, 16'd53CC, 16'd32C8, 16'd11C5, 16'd0102, 16'd00A0, 16'd0060, 16'd0060, 16'd0040, 16'd0040, 16'd0040, 16'd0060, 16'd0080, 16'd0080, 16'd0081, 16'd0081, 16'd0081, 16'd0061, 16'd0040, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0861, 16'd1964, 16'd3268, 16'd4B4B, 16'd53CD, 16'd53CD, 16'd53AC, 16'd4B8B, 16'd4B6B, 16'd4B6B, 16'd4B8B, 16'd4B8B, 16'd4B4B, 16'd3AC8, 16'd2206, 16'd0963, 16'd00E1, 16'd0080, 16'd0060, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0060, 16'd0060, 16'd0060, 16'd0060, 16'd0060, 16'd0040, 16'd0040, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0040, 16'd10E2, 16'd1985, 16'd2A26, 16'd2A67, 16'd2A67, 16'd2A27, 16'd2A06, 16'd2A06, 16'd2A06, 16'd2A26, 16'd2A26, 16'd2206, 16'd19A5, 16'd1143, 16'd00E2, 16'd00A0, 16'd0060, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0061, 16'd08C2, 16'd0902, 16'd0923, 16'd0923, 16'd0902, 16'd08E2, 16'd08E1, 16'd08E1, 16'd08E2, 16'd08E2, 16'd08E2, 16'd08C1, 16'd00A1, 16'd0080, 16'd0060, 16'd0060, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0040, 16'd0060, 16'd0060, 16'd0060, 16'd0040, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0040, 16'd0060, 16'd0861, 16'd0861, 16'd0040, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0040, 16'd0861, 16'd0881, 16'd0881, 16'd0860, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0040, 16'd0881, 16'd0881, 16'd0881, 16'd0861, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0060, 16'd0861, 16'd0881, 16'd0861, 16'd0040, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0820, 16'd0840, 16'd0841, 16'd0840, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0040, 16'd0840, 16'd0840, 16'd0860, 16'd0861, 16'd0860, 16'd0040, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0841, 16'd1061, 16'd1061, 16'd0861, 16'd0820, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0840, 16'd0861, 16'd0861, 16'd0861, 16'd0860, 16'd0040, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0840, 16'd1061, 16'd1081, 16'd1082, 16'd1061, 16'd0840, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0840, 16'd0860, 16'd0861, 16'd0881, 16'd0881, 16'd0860, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0840, 16'd1061, 16'd1082, 16'd18A2, 16'd1081, 16'd0840, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0840, 16'd0860, 16'd0881, 16'd1081, 16'd0881, 16'd0840, 16'd0020, 16'd0000, 16'd0020, 16'd0040, 16'd0061, 16'd0881, 16'd0881, 16'd0061, 16'd0040, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0820, 16'd0861, 16'd1081, 16'd1081, 16'd1061, 16'd0840, 16'd0820, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0840, 16'd0861, 16'd0881, 16'd0861, 16'd0040, 16'd0000, 16'd0000, 16'd0040, 16'd10A2, 16'd1924, 16'd2165, 16'd2164, 16'd1903, 16'd08A1, 16'd0040, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0841, 16'd1061, 16'd1061, 16'd0841, 16'd0820, 16'd0820, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0820, 16'd0840, 16'd0861, 16'd0840, 16'd0020, 16'd0000, 16'd0020, 16'd0881, 16'd2144, 16'd3A27, 16'd4A89, 16'd4269, 16'd31E6, 16'd1903, 16'd0060, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0820, 16'd0820, 16'd0820, 16'd0820, 16'd0820, 16'd0820, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0020, 16'd10E2, 16'd3207, 16'd5B2B, 16'd73CE, 16'd6BAD, 16'd4AAA, 16'd2965, 16'd0861, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0820, 16'd0820, 16'd0820, 16'd0820, 16'd0820, 16'd0820, 16'd0820, 16'd0820, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0040, 16'd1923, 16'd4AA9, 16'd740F, 16'd94F2, 16'd8CB1, 16'd636D, 16'd31E6, 16'd0881, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0820, 16'd0820, 16'd0820, 16'd0820, 16'd0820, 16'd0820, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0040, 16'd1944, 16'd530B, 16'd8CB1, 16'dADB5, 16'dA574, 16'd73EF, 16'd3A27, 16'd0881, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0820, 16'd0820, 16'd0820, 16'd0820, 16'd0800, 16'd0820, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0040, 16'd2164, 16'd5B2B, 16'd9513, 16'dB617, 16'dADD6, 16'd7C50, 16'd4248, 16'd08A1, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd2164, 16'd5B4C, 16'd9D33, 16'dBE58, 16'dB5F7, 16'd8470, 16'd4248, 16'd08A1, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd2144, 16'd5B4C, 16'd9D33, 16'dBE58, 16'dB617, 16'd8471, 16'd4268, 16'd08A1, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd2144, 16'd5B2B, 16'd9533, 16'dBE58, 16'dB617, 16'd8470, 16'd4268, 16'd08A1, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0040, 16'd0060, 16'd0060, 16'd0060, 16'd0040, 16'd0040, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd1924, 16'd5B2B, 16'd9533, 16'dBE58, 16'dB617, 16'd8470, 16'd4268, 16'd08A1, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0060, 16'd0060, 16'd0060, 16'd0060, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd1923, 16'd5B2B, 16'd9513, 16'dB657, 16'dADF6, 16'd7C70, 16'd4268, 16'd08A1, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0060, 16'd0060, 16'd0060, 16'd0040, 16'd0000, 16'd0000, 16'd0000, 16'd1923, 16'd530B, 16'd8CF2, 16'dB617, 16'dA5D6, 16'd7C50, 16'd3A48, 16'd08A1, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0060, 16'd0060, 16'd0040, 16'd0000, 16'd0000, 16'd0020, 16'd1923, 16'd52EA, 16'd8CD2, 16'dADF6, 16'dA595, 16'd742F, 16'd3A48, 16'd08A1, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0060, 16'd0060, 16'd0040, 16'd0000, 16'd0000, 16'd0020, 16'd1923, 16'd4AEA, 16'd84B1, 16'dA5B5, 16'd9D74, 16'd740F, 16'd3A27, 16'd08A1, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0060, 16'd0080, 16'd0060, 16'd0000, 16'd0000, 16'd0020, 16'd1923, 16'd4ACA, 16'd8491, 16'd9D95, 16'd9554, 16'd6BEE, 16'd3A27, 16'd08A1, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0000, 16'd0020, 16'd0040, 16'd0060, 16'd0080, 16'd0060, 16'd0000, 16'd0000, 16'd0020, 16'd1923, 16'd4ACA, 16'd7C90, 16'd9D95, 16'd9553, 16'd6BEE, 16'd3A27, 16'd08A1, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0000, 16'd0000, 16'd0020, 16'd0040, 16'd0060, 16'd0080, 16'd0060, 16'd0000, 16'd0000, 16'd0020, 16'd1923, 16'd4ACA, 16'd7C90, 16'd9D94, 16'd9533, 16'd6BEE, 16'd3A27, 16'd08A1, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0000, 16'd0000, 16'd0020, 16'd0040, 16'd0060, 16'd0080, 16'd0060, 16'd0000, 16'd0000, 16'd0020, 16'd1923, 16'd4ACA, 16'd7C90, 16'd9D94, 16'd9533, 16'd6BEE, 16'd3A27, 16'd08A1, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0000, 16'd0020, 16'd0040, 16'd0060, 16'd0080, 16'd0060, 16'd0000, 16'd0000, 16'd0020, 16'd1923, 16'd4ACA, 16'd7C90, 16'd9D95, 16'd9553, 16'd6BEE, 16'd3A27, 16'd08A1, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0060, 16'd0080, 16'd0060, 16'd0000, 16'd0000, 16'd0020, 16'd1923, 16'd4ACA, 16'd8491, 16'd9D95, 16'd9554, 16'd6BEE, 16'd3A27, 16'd08A1, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0060, 16'd0060, 16'd0040, 16'd0000, 16'd0000, 16'd0020, 16'd1923, 16'd4AEA, 16'd84B1, 16'dA5B5, 16'd9D74, 16'd740F, 16'd3A27, 16'd08A1, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0060, 16'd0060, 16'd0040, 16'd0000, 16'd0000, 16'd0020, 16'd1923, 16'd52EA, 16'd8CD2, 16'dADF6, 16'dA595, 16'd742F, 16'd3A48, 16'd08A1, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0060, 16'd0060, 16'd0060, 16'd0040, 16'd0000, 16'd0000, 16'd0000, 16'd1923, 16'd530B, 16'd8CF2, 16'dB617, 16'dA5D6, 16'd7C50, 16'd3A48, 16'd08A1, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0060, 16'd0060, 16'd0060, 16'd0060, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd1923, 16'd5B2B, 16'd9513, 16'dB657, 16'dADF6, 16'd7C70, 16'd4268, 16'd08A1, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0040, 16'd0060, 16'd0060, 16'd0060, 16'd0040, 16'd0040, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd1924, 16'd5B2B, 16'd9533, 16'dBE58, 16'dB617, 16'd8470, 16'd4268, 16'd08A1, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd2144, 16'd5B2B, 16'd9533, 16'dBE58, 16'dB617, 16'd8470, 16'd4268, 16'd08A1, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd2144, 16'd5B4C, 16'd9D33, 16'dBE58, 16'dB617, 16'd8471, 16'd4268, 16'd08A1, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd2164, 16'd5B4C, 16'd9D33, 16'dBE58, 16'dB5F7, 16'd8470, 16'd4248, 16'd08A1, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0820, 16'd0820, 16'd0820, 16'd0820, 16'd0800, 16'd0820, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0040, 16'd2164, 16'd5B2B, 16'd9513, 16'dB617, 16'dADD6, 16'd7C50, 16'd4248, 16'd08A1, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0820, 16'd0820, 16'd0820, 16'd0820, 16'd0820, 16'd0820, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0040, 16'd1944, 16'd530B, 16'd8CB1, 16'dADB5, 16'dA574, 16'd73EF, 16'd3A27, 16'd0881, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0820, 16'd0820, 16'd0820, 16'd0820, 16'd0820, 16'd0820, 16'd0820, 16'd0820, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0040, 16'd1923, 16'd4AA9, 16'd740F, 16'd94F2, 16'd8CB1, 16'd636D, 16'd31E6, 16'd0881, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0820, 16'd0820, 16'd0820, 16'd0820, 16'd0820, 16'd0820, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0020, 16'd10E2, 16'd3207, 16'd5B2B, 16'd73CE, 16'd6BAD, 16'd4AAA, 16'd2965, 16'd0861, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0841, 16'd1061, 16'd1061, 16'd0841, 16'd0820, 16'd0820, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0820, 16'd0840, 16'd0861, 16'd0840, 16'd0020, 16'd0000, 16'd0020, 16'd0881, 16'd2144, 16'd3A27, 16'd4A89, 16'd4269, 16'd31E6, 16'd1903, 16'd0060, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0820, 16'd0861, 16'd1081, 16'd1081, 16'd1061, 16'd0840, 16'd0820, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0840, 16'd0861, 16'd0881, 16'd0861, 16'd0040, 16'd0000, 16'd0000, 16'd0040, 16'd10A2, 16'd1924, 16'd2165, 16'd2164, 16'd1903, 16'd08A1, 16'd0040, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0840, 16'd1061, 16'd1082, 16'd18A2, 16'd1081, 16'd0840, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0840, 16'd0860, 16'd0881, 16'd1081, 16'd0881, 16'd0840, 16'd0020, 16'd0000, 16'd0020, 16'd0040, 16'd0061, 16'd0881, 16'd0881, 16'd0061, 16'd0040, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0840, 16'd1061, 16'd1081, 16'd1082, 16'd1061, 16'd0840, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0840, 16'd0860, 16'd0861, 16'd0881, 16'd0881, 16'd0860, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0841, 16'd1061, 16'd1061, 16'd0861, 16'd0820, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0840, 16'd0861, 16'd0861, 16'd0861, 16'd0860, 16'd0040, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0820, 16'd0840, 16'd0841, 16'd0840, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0040, 16'd0840, 16'd0840, 16'd0860, 16'd0861, 16'd0860, 16'd0040, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0060, 16'd0861, 16'd0881, 16'd0861, 16'd0040, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0040, 16'd0881, 16'd0881, 16'd0881, 16'd0861, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0040, 16'd0861, 16'd0881, 16'd0881, 16'd0860, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0040, 16'd0060, 16'd0861, 16'd0861, 16'd0040, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0040, 16'd0060, 16'd0060, 16'd0060, 16'd0040, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0061, 16'd08C2, 16'd0902, 16'd0923, 16'd0923, 16'd0902, 16'd08E2, 16'd08E1, 16'd08E1, 16'd08E2, 16'd08E2, 16'd08E2, 16'd08C1, 16'd00A1, 16'd0080, 16'd0060, 16'd0060, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0040, 16'd10E2, 16'd1985, 16'd2A26, 16'd2A67, 16'd2A67, 16'd2A27, 16'd2A06, 16'd2A06, 16'd2A06, 16'd2A26, 16'd2A26, 16'd2206, 16'd19A5, 16'd1143, 16'd00E2, 16'd00A0, 16'd0060, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0861, 16'd1964, 16'd3268, 16'd4B4B, 16'd53CD, 16'd53CD, 16'd53AC, 16'd4B8B, 16'd4B6B, 16'd4B6B, 16'd4B8B, 16'd4B8B, 16'd4B4B, 16'd3AC8, 16'd2206, 16'd0963, 16'd00E1, 16'd0080, 16'd0060, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0060, 16'd0060, 16'd0060, 16'd0060, 16'd0060, 16'd0040, 16'd0040, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0881, 16'd29C6, 16'd534B, 16'd6C90, 16'd7D32, 16'd7D52, 16'd7511, 16'd6CF0, 16'd6CD0, 16'd6CD0, 16'd74F1, 16'd74D1, 16'd6C8F, 16'd53CC, 16'd32C8, 16'd11C5, 16'd0102, 16'd00A0, 16'd0060, 16'd0060, 16'd0040, 16'd0040, 16'd0040, 16'd0060, 16'd0080, 16'd0080, 16'd0081, 16'd0081, 16'd0081, 16'd0061, 16'd0040, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd08A2, 16'd3247, 16'd640E, 16'd8D94, 16'd9E56, 16'd9E77, 16'd9636, 16'd8DF4, 16'd85D4, 16'd8DF4, 16'd8E15, 16'd8DF5, 16'd8593, 16'd648F, 16'd3B4B, 16'd1A06, 16'd0122, 16'd00A0, 16'd0080, 16'd0060, 16'd0040, 16'd0040, 16'd0060, 16'd0080, 16'd0081, 16'd00A1, 16'd00A1, 16'd00A1, 16'd00A1, 16'd0081, 16'd0061, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd10C2, 16'd3A88, 16'd7490, 16'd9E36, 16'dB719, 16'dB739, 16'dA6F8, 16'd9E97, 16'd9676, 16'd9E97, 16'd9EB7, 16'd9EB7, 16'd9636, 16'd7511, 16'd43AC, 16'd1A26, 16'd0122, 16'd00A0, 16'd0060, 16'd0060, 16'd0060, 16'd0060, 16'd0060, 16'd0080, 16'd00A1, 16'd00A1, 16'd00A1, 16'd00A1, 16'd0081, 16'd0081, 16'd0061, 16'd0040, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd10E2, 16'd42A9, 16'd7CF1, 16'dAEB8, 16'dBF9B, 16'dBFBB, 16'dAF59, 16'd9ED8, 16'd96B7, 16'd9ED8, 16'dA718, 16'dA719, 16'd9E97, 16'd7D52, 16'd4BAC, 16'd1A26, 16'd0102, 16'd0080, 16'd0060, 16'd0060, 16'd0060, 16'd0060, 16'd0060, 16'd0080, 16'd00A0, 16'd00A0, 16'd0081, 16'd0081, 16'd0081, 16'd0061, 16'd0061, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd10E2, 16'd42EA, 16'd8512, 16'dB719, 16'dC7DC, 16'dC7DC, 16'dAF7A, 16'd9EF8, 16'd96B7, 16'd9EF8, 16'dA739, 16'dAF39, 16'd9EB7, 16'd7D73, 16'd4BAC, 16'd1A05, 16'd00E1, 16'd0060, 16'd0040, 16'd0060, 16'd0060, 16'd0060, 16'd0080, 16'd0080, 16'd0080, 16'd0080, 16'd0060, 16'd0060, 16'd0060, 16'd0040, 16'd0040, 16'd0061, 16'd0861, 16'd0841, 16'd0040, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd10E2, 16'd4AEA, 16'd8553, 16'dB73A, 16'dCFFD, 16'dC7FC, 16'dAF7A, 16'd9ED7, 16'd96B6, 16'd96D7, 16'dA739, 16'dAF59, 16'd9ED8, 16'd7D73, 16'd4BAC, 16'd19E5, 16'd00A0, 16'd0040, 16'd0040, 16'd0060, 16'd0080, 16'd0080, 16'd0080, 16'd0080, 16'd0080, 16'd0060, 16'd0060, 16'd0040, 16'd0020, 16'd0040, 16'd0040, 16'd0861, 16'd0881, 16'd0881, 16'd0841, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd10E2, 16'd4B0A, 16'd8553, 16'dB75A, 16'dCFFD, 16'dC7FC, 16'dAF7A, 16'd96D7, 16'd8E96, 16'd96D7, 16'dA739, 16'dA759, 16'd9ED8, 16'd7D72, 16'd4B8B, 16'd19C4, 16'd0080, 16'd0020, 16'd0020, 16'd0060, 16'd0080, 16'd0080, 16'd0080, 16'd0080, 16'd0060, 16'd0060, 16'd0040, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0881, 16'd08A2, 16'd0881, 16'd0861, 16'd0840, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd10E2, 16'd4B0A, 16'd8553, 16'dB75A, 16'dCFFD, 16'dC7FC, 16'dAF7A, 16'd96D7, 16'd8E96, 16'd96D7, 16'dA739, 16'dA75A, 16'd9ED8, 16'd7D72, 16'd4B8B, 16'd19A4, 16'd0080, 16'd0020, 16'd0020, 16'd0060, 16'd0080, 16'd0080, 16'd0080, 16'd0060, 16'd0060, 16'd0060, 16'd0040, 16'd0020, 16'd0020, 16'd0040, 16'd0061, 16'd0881, 16'd08A2, 16'd0881, 16'd0861, 16'd0840, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd10E2, 16'd42EA, 16'd8553, 16'dB73A, 16'dC7FD, 16'dC7FC, 16'dAF9A, 16'd96F8, 16'd8ED7, 16'd96F8, 16'dA759, 16'dAF7A, 16'd9ED8, 16'd7D72, 16'd4B8B, 16'd19C4, 16'd0080, 16'd0020, 16'd0020, 16'd0060, 16'd0080, 16'd0080, 16'd0080, 16'd0060, 16'd0060, 16'd0060, 16'd0040, 16'd0040, 16'd0060, 16'd0061, 16'd0861, 16'd0881, 16'd0881, 16'd0861, 16'd0841, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd10E2, 16'd42E9, 16'd7D32, 16'dAF19, 16'dC7FC, 16'dBFFC, 16'dAF9A, 16'd9F18, 16'd96F7, 16'd9F38, 16'dA759, 16'dA77A, 16'd9ED8, 16'd7D72, 16'd4BAB, 16'd19C4, 16'd00A0, 16'd0020, 16'd0020, 16'd0060, 16'd0080, 16'd0080, 16'd0060, 16'd0060, 16'd0040, 16'd0060, 16'd0060, 16'd0881, 16'd08A1, 16'd08A1, 16'd0881, 16'd0861, 16'd0861, 16'd0841, 16'd0040, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd10E2, 16'd42C9, 16'd74F1, 16'dA6D8, 16'dB7BB, 16'dB7DB, 16'dAF9A, 16'd9F38, 16'd96F8, 16'd9F38, 16'dA759, 16'dA759, 16'd96B7, 16'd7572, 16'd4B8B, 16'd19E4, 16'd00C0, 16'd0040, 16'd0040, 16'd0060, 16'd0080, 16'd0060, 16'd0060, 16'd0040, 16'd0040, 16'd0060, 16'd0881, 16'd08C2, 16'd10E2, 16'd10C2, 16'd08A2, 16'd0861, 16'd0040, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd10C2, 16'd3A88, 16'd6C90, 16'd9656, 16'dAF39, 16'dAF5A, 16'dA739, 16'd96F7, 16'd96D7, 16'd96F8, 16'd9F18, 16'd9EF8, 16'd8E76, 16'd6D31, 16'd438B, 16'd19E4, 16'd00C0, 16'd0040, 16'd0040, 16'd0060, 16'd0080, 16'd0060, 16'd0060, 16'd0040, 16'd0040, 16'd0060, 16'd08A1, 16'd10C2, 16'd1103, 16'd10E3, 16'd08A2, 16'd0861, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd08C2, 16'd3247, 16'd5C0E, 16'd8593, 16'd9676, 16'd9697, 16'd8E76, 16'd8655, 16'd8635, 16'd8655, 16'd8E76, 16'd8E56, 16'd7DD4, 16'd64AF, 16'd3B29, 16'd11C4, 16'd00C0, 16'd0060, 16'd0040, 16'd0060, 16'd0080, 16'd0060, 16'd0040, 16'd0040, 16'd0040, 16'd0060, 16'd0881, 16'd10C2, 16'd1103, 16'd10E3, 16'd08A2, 16'd0041, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd08A1, 16'd29E6, 16'd4B4B, 16'd648F, 16'd7531, 16'd7552, 16'd7551, 16'd6D31, 16'd6D10, 16'd6D51, 16'd6D52, 16'd6D52, 16'd64F0, 16'd4C0D, 16'd2AC8, 16'd1183, 16'd00C0, 16'd0060, 16'd0040, 16'd0060, 16'd0060, 16'd0060, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0881, 16'd08A2, 16'd10C2, 16'd10C2, 16'd0881, 16'd0040, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0081, 16'd1964, 16'd3267, 16'd432A, 16'd4BAC, 16'd53CC, 16'd4BCC, 16'd4BAB, 16'd43AB, 16'd4BEC, 16'd4C0D, 16'd4C0D, 16'd43CC, 16'd3329, 16'd2226, 16'd0942, 16'd00A0, 16'd0040, 16'd0040, 16'd0060, 16'd0060, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0040, 16'd0060, 16'd0881, 16'd08A2, 16'd0881, 16'd0861, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0040, 16'd08E2, 16'd1964, 16'd21E5, 16'd2A46, 16'd2A46, 16'd2A46, 16'd2246, 16'd2246, 16'd2287, 16'd2AA8, 16'd2AC8, 16'd22C8, 16'd1A46, 16'd11A4, 16'd00E1, 16'd0080, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0061, 16'd0041, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0040, 16'd0060, 16'd08A1, 16'd08E1, 16'd0901, 16'd0901, 16'd0901, 16'd0901, 16'd0921, 16'd0942, 16'd0983, 16'd09C4, 16'd09C4, 16'd0983, 16'd0122, 16'd00A0, 16'd0060, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0060, 16'd00A0, 16'd00E1, 16'd0101, 16'd0122, 16'd0101, 16'd00C1, 16'd0080, 16'd0060, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0040, 16'd0080, 16'd00A0, 16'd00C0, 16'd00C0, 16'd00A0, 16'd0080, 16'd0060, 16'd0060, 16'd0060, 16'd0060, 16'd0060, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0040, 16'd0060, 16'd0080, 16'd0080, 16'd0080, 16'd0080, 16'd0080, 16'd0080, 16'd0080, 16'd0080, 16'd0060, 16'd0060, 16'd0060, 16'd0060, 16'd0060, 16'd0040, 16'd0040, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0060, 16'd0060, 16'd0080, 16'd0080, 16'd0080, 16'd0080, 16'd0080, 16'd0081, 16'd0081, 16'd0081, 16'd0081, 16'd0080, 16'd0060, 16'd0060, 16'd0040, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0840, 16'd0840, 16'd0820, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0060, 16'd0060, 16'd0060, 16'd0080, 16'd0080, 16'd0081, 16'd00A1, 16'd00A1, 16'd00A1, 16'd0081, 16'd0081, 16'd0081, 16'd0081, 16'd0060, 16'd0040, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0840, 16'd0841, 16'd0841, 16'd0840, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0060, 16'd0080, 16'd0081, 16'd00A1, 16'd00A1, 16'd00A1, 16'd0081, 16'd0081, 16'd0081, 16'd0081, 16'd0060, 16'd0040, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0840, 16'd0841, 16'd0841, 16'd0840, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0060, 16'd0080, 16'd0081, 16'd0081, 16'd0081, 16'd0081, 16'd0061, 16'd0061, 16'd0060, 16'd0040, 16'd0040, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0820, 16'd0841, 16'd0841, 16'd0820, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0060, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0060, 16'd0060, 16'd0060, 16'd0060, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0820, 16'd0820, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0040, 16'd0040, 16'd0060, 16'd0060, 16'd0060, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0040,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0040, 16'd0060, 16'd0060, 16'd0060, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0040,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0040, 16'd0060, 16'd0060, 16'd0060, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0040,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0040,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0820, 16'd0800, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0040,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0820, 16'd0820, 16'd0820, 16'd0820, 16'd0820, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0040,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0820, 16'd0820, 16'd0820, 16'd0841, 16'd0821, 16'd0820, 16'd0800, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0820, 16'd0820, 16'd0820, 16'd0841, 16'd0821, 16'd0820, 16'd0800, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0820, 16'd0820, 16'd0820, 16'd0820, 16'd0800, 16'd0800, 16'd0800, 16'd0820, 16'd0820, 16'd0820, 16'd0820, 16'd0820, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0820, 16'd0820, 16'd0840, 16'd0820, 16'd0820, 16'd0820, 16'd0000, 16'd0000, 16'd0820, 16'd0820, 16'd0820, 16'd0820, 16'd0800, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0820, 16'd0820, 16'd0840, 16'd0840, 16'd0840, 16'd0820, 16'd0820, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0820, 16'd0820, 16'd1041, 16'd1061, 16'd0841, 16'd0840, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0820, 16'd0840, 16'd1061, 16'd1061, 16'd0841, 16'd0840, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0820, 16'd0840, 16'd0861, 16'd1061, 16'd0841, 16'd0840, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0840, 16'd0861, 16'd0861, 16'd0841, 16'd0840, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0840, 16'd0840, 16'd0861, 16'd0840, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0840, 16'd0840, 16'd0840, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0040, 16'd0840, 16'd0040, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0840, 16'd0840, 16'd0820, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0840, 16'd0840, 16'd0820, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0040, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0840, 16'd0840, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0040, 16'd0840, 16'd0840, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0040, 16'd0060, 16'd0060, 16'd0060, 16'd0040, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0040, 16'd0060, 16'd0060, 16'd0080, 16'd0060, 16'd0040, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0040, 16'd0060, 16'd0081, 16'd0081, 16'd0060, 16'd0040, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000,
        16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0040, 16'd0060, 16'd0081, 16'd0081, 16'd0060, 16'd0040, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0020, 16'd0020, 16'd0020, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0020, 16'd0040, 16'd0040, 16'd0040, 16'd0020, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0000, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd0800, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000, 16'd1000,
    };
    reg [0:15] img_out [21384:0];

    always @(*) begin
        if(step == 0) img_out <= step0;
        else img_out <= img_out;
    end

    assign ram_data = img_out[ram_addr_y*132 + ram_addr_x];
    
endmodule