module smile (
    input wire clk,
    input wire rst,
    input wire [7:0] ram_addr,
    output wire [131:0] ram_data
);

    
    
endmodule